module leds_alarm (Y, led_a, led_b, led_c, led_d, led_e, led_f, led_g, led_h, led_i, led_j);
  input Y;
  output led_a, led_b, led_c, led_d, led_e, led_f, led_g, led_h, led_i, led_j;
  
   assign led_a = Y;
   assign led_b = Y;
   assign led_c = Y;
   assign led_d = Y;
   assign led_e = Y;
   assign led_f = Y;
   assign led_g = Y;
   assign led_h = Y;
   assign led_i = Y;
   assign led_j = Y;
  
endmodule